// Параметрическое задание разрядности счетчика
`define m 4

// Схема суммирующего декадного счетчика с синхронным сбросом в ноль 
// и с входом 'ce' разрешения счета
module VCDmRE (

  input ce,  // Clock Enable - сигнал разрешения счета
  input clk, // Сигнал синхронизации (тактирующий сигнал)
  input R,   // Сигнал синхронного сброса в ноль

  output reg [`m-1:0]Q = 0, // Значение счетчика
  output wire TC,           // Terminal Count - сигнал переполнения
  output wire CEO           // Clock Enable Output - сигнал переноса
);

// Q0 & Q1 &...& Q'm-1 == 1
assign TC = (Q == 9);

// Сигнал переноса
assign CEO = ce & TC;

// По фронту входа синхронизации
always @(posedge clk) begin
  
  // Сброс в 0 происходит при при Q == 9 и ce == 1 или при R == 1
  // Иначе если ce == 1, то "суммировать", иначе "стоять"
  Q <= (R | CEO)? 0 : ce? Q+1 : Q;
end

endmodule
