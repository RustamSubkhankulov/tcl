`timescale 1ns / 1ps

module MASTER_I2C(

  inout SDA,                     // Физический сигнал 'SDA' мастера
  input st,                      // Импульс запуска передачи
  input clk,                     // Сигнал синхронизации
  
  input [7:0]ADR_COM,            // Адрес-команда (адрес ведомого + команда)
                                 // [7:1] - адрес ведомого
                                 // [0] - команда: 0 - запись, 1 - чтение

  input [7:0]adr_REG,            // Адрес регистра ведомого
  input [7:0]dat_REG,            // Данные для ведомого


  output reg SCL            = 1, // Сигнал SCL мастера
  output reg SDA_MASTER     = 1, // Логический сигнал 'SDA' мастера
  
  output reg T_start        = 0, // Старт передачи
  output reg T_stop         = 0, // Стоп передачи
  
  output reg [3:0]cb_bit    = 0, // Счетчик бит
  output reg en_tx          = 0, // Разрешение передачи
  
  output wire ce_tact,           // Границы тактов
  output wire ce_bit,            // Середины тактов
  output wire ce_byte,           // Границы байт

  output wire T_AC,              // Такт подтверждения  
  output wire ce_AC,             // Строб такта 'T_AC'
  output wire err_AC,            // Триггер подтверждения
  
  output reg [2:0]cb_byte   = 0, // Счетчик байт
  
  output reg [7:0]sr_rx_SDA = 0, // Регистр сдвига принимаемых данных
  output reg [7:0]RX_dat    = 0  // Регистр данных от ведомого
);

// PULLUP Резистор
PULLUP DA1(SDA);

// Выходной буфер с третьим состоянием (SDA=SDA_MASTER & SDA_SLAVE)
BUFT DD1(.I(1'b0), .O(SDA), .T(SDA_MASTER))

parameter Fclk   = 50000000;          // Fclk = 50000 kHz
parameter Fvel   = 1250000;           // Fvel = 1250 kHz
parameter N4vel  = Fclk / (4 * Fvel); // 50000000 / (4 * 1250000) = 10
parameter N_byte = 3 ;                // Число байт (адрес ведомого, адрес регистра, данные)

reg [10:0]cb_ce = 4 * N4vel;
assign ce_tact  = (cb_ce == 1 * N4vel);         // 10, границы тактов
assign ce_bit   = (cb_ce == 3 * N4vel) & en_tx; // 30, середины тактов

reg [7:0]sr_tx_SDA = 8'h00 ; // Регистр сдвига передаваемых данных

assign T_AC  = (cb_bit == 8);                      // Такт подтверждения
wire   T_dat = en_tx & !T_start & !T_stop & !T_AC; // Такт передачи данных

assign ce_AC   = T_AC & ce_bit;                    // Строб такта 'T_AC'
assign ce_byte = ce_tact & T_AC;                   // Границы байт

wire R_W = ADR_COM[0]; // Команда: 1-чтение, 0-запись
reg rep_st = 0;        // ?

wire [7:0]TX_dat = (cb_byte == 0)?          ADR_COM : // Адрес-команда
                   (cb_byte == 1)?          adr_REG : // Адрес регистра
                   ((cb_byte == 2) & !R_W)? dat_REG : // Данные регистра
                   8'hFF ; 

always @ (posedge clk) begin
  
  // 3 * N4vel - задержка первого (следующего) 'ce_bit' от 'st'
  // При импульсе запуска передачи устанавливаем задержку первого 'ce_bit'.
  // Если значение счетчика дошло до 0, устанавливаем 4 * N4vel,
  // иначе декрементируем значение счетчика по сигналу синхронизации.
  cb_ce <= st? 3 * N4vel : (cb_ce == 1)? 4 * N4vel : cb_ce-1 ; 
  
  // Старт передачи (уст. в единицу) при импульсе запуска передачи, 
  // иначе по границе такта устанавливаем в ноль (такт не является тактом старта передачи)
  T_start <= st? 1 : ce_tact? 0 : T_start;
  
  // Сбрасываем счётчик битов в 0 при импульсе запуска передачи или по границе байта.
  // Иначе по границе такта (кроме стартового) при разрешенной передаче инкрементируем.
  cb_bit <= (st | ce_byte)? 0 : (ce_tact & en_tx & !T_start)? cb_bit+1 : cb_bit;
  
  // Стоп передачи при: граница байта, при этом байт последний в кадре
  // или не было получено подтверждение от ведомого.
  // Иначе по стробу такта выставляем в ноль (передача продолжается)
  T_stop <= ce_byte & ((cb_byte == N_byte - 1) | err_AC)? 1 : ce_bit? 0 : T_stop;
  
  // Разрешение передачи выставляем по импульсу запуска передачи,
  // Выставялем в ноль в случае завершения передачи по стробу такта.
  en_tx <= st? 1 : (T_stop & ce_bit)? 0 : en_tx;
  
  // Сигнал синхронизации высокий при запрещенной передаче
  // При разрешенной передаче высокий в промежутке (2 * N4vel; 1] счетчика 'cb_ce'.
  SCL <= (cb_ce > 2*N4vel) | !en_tx;

  // Устанавливаем 0 при старте передачи или перед завершением.
  // Иначе при разрешенной передаче на тактах передачи данных выставляем
  // бит данных из сдвигового регистра, на такте подтверждения - единицу.
  // Иначе линия установлена в единицу.
  SDA_MASTER <= (T_start | T_stop)? 0 : en_tx? (sr_tx_SDA[7] | T_AC) : 1;
  
  // Загружаем данные в сдвиговый регистр по необходимости, 
  // иначе производим непосредственно сдвиг данных в регистре.
  sr_tx_SDA <= rep_st? TX_dat : (ce_tact & T_dat)? sr_tx_SDA<<1 | 1'b1 : sr_tx_SDA;
  
  // Обновляем значение счётчика байтов.
  cb_byte <= st? 0 : (ce_byte & en_tx)? cb_byte+1 : cb_byte;
  
  // Триггер подтверждения сбрасывается по имппульсу запуска передачи
  // По стробу такта подтверждения, если ведомый не отправил подтверждение,
  // устанавливаем в 1 - нет подтверждения.
  err_AC <= st? 0 : (ce_AC & SDA)? 1 : err_AC;
  
  // Сигнал загрузки данных для отправки, устанавливается по импульсу запуска
  // передачи, или при отправке следующего байта данных при условии, что передача
  // разерешена.
  rep_st = (st | (ce_byte & en_tx));
  
  // Последовательный прием данных от ведомого на интервале третьего байта
  sr_rx_SDA <= ((cb_byte == N_byte-1) & ce_bit & T_dat)? sr_rx_SDA<<1 | SDA : sr_rx_SDA;

  // Загружаем данные от ведомого по завершении третьего байта при команде 'чтение'
  RX_dat <= ((cb_byte == N_byte-1) & ce_byte & R_W)? sr_rx_SDA : RX_dat;
end

endmodule // MASTER_I2C