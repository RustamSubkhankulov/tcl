// Параметрическое задание разрядности счетчика
`define m 4

// Схема m-разрядного реверсивного счетчика с асинхронным сбросом в ноль
module VCBmCLED (

  input ce,          // Clock Enable - сигнал разрешения счета
  input up,          // Направление счета
  input [`m-1:0] di, // Значение счетчика при загрузке
  input L,           // Сигнал разрешения синхронной загрузки
  input clk,         // Сигнал синхронизации (тактирующий сигнал)
  input clr,         // Сигнал асинхронного сброса в ноль

  output reg [`m-1:0] Q = 0, // Значение счетчика
  output wire TC,            // Terminal Count - сигнал переполнения
  output wire CEO            // Clock Enable Output - сигнал переноса
);

// Q0 & Q1 &...& Q'm-1 == 1 при up == 1
// Q0 & Q1 &...& Q'm-1 == 0 при up == 0
assign TC = up? (Q == ((1 << `m) - 1)) : (Q == 0);

// Сигнал переноса
assign CEO = ce & TC;

// По фронту входа синхронизации или по фронту сигнала асинхронного сброса
always @ (posedge clr or posedge clk) begin
  
  // Асинхронный сброс
  if (clr) Q <= 0;
  // При clr == L == 0, ce == 1, up == 1 "суммировать"
  // При clr == L == 0, ce == 1, up == 0 "вычитать"
  // При clr == 0, L == 1 независимо от ce значение  счетчика выставляется в di
  else     Q <= L? di : (up & ce)? Q+1 : (!up & ce)? Q-1 : Q; 
end

endmodule
