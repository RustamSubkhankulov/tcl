// Параметрическое задание разрядности счетчика
`define m 4

// Схема m-разрядного счетчика Джонсона с синхронным сбросом в ноль 
// и с входом 'ce' разрешения счета
module VCJmRE (

  input ce,  // Clock Enable - сигнал разрешения счета
  input clk, // Сигнал синхронизации (тактирующий сигнал)
  input R,   // Сигнал синхронного сброса в ноль

  output reg [`m-1:0] Q = 0, // Значение счетчика
  output wire TC,            // Terminal Count - сигнал переполнения
  output wire CEO            // Clock Enable Output - сигнал переноса
);

// Q0 & Q1 &...& Q'm-1 == 1
assign TC = (Q == (1 << `m) - 1);

// Сигнал переноса
assign CEO = ce & TC;

// По фронту входа синхронизации
always @ (posedge clk) begin
  
  // Если R == 1, то сброс в 0 независимо от сигнала синхронизации clk
  // Иначе переходим к следующей итерации цикла 
  // (в счетчике Джонсона возможно несколько устойчивых циклов)
  Q <= R? 0 : ce? (Q << 1) | (!Q[`m-1]) : Q;
end

endmodule
