// Параметрическое задание разрядности счетчика
`define m 4

// Схема вычитающего m-разрядного счетчика с синхронным сбросом в ноль 
// и с входом 'ce' разрешения счета
module VCBDmSE (

  input ce,  // Clock Enable - сигнал разрешения счета
  input clk, // Сигнал синхронизации (тактирующий сигнал)
  input s,   // Сигнал синхронной установки в 2^m-1

  output reg [`m-1:0]Q = 0, // Значение счетчика
  output wire TC,           // Terminal Count - сигнал переполнения
  output wire CEO           // Clock Enable Output - сигнал переноса
);

// Q0 & Q1 &...& Q'm-1 == 0
assign TC = (Q == 0);

// Сигнал переноса
assign CEO = ce & TC;

// По фронту входа синхронизации
always @(posedge clk) begin
  
  // Если s == 1, то запись 2^m-1
  // Иначе если ce == 1, то "вычитать", иначе "стоять"
  Q <= (s)? ((1 << `m) - 1) : ce? Q-1 : Q;
end

endmodule
